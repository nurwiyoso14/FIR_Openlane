VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO shifter
  CLASS BLOCK ;
  FOREIGN shifter ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 789.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 796.000 398.520 800.000 399.120 ;
    END
  END clk
  PIN input_pc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 27.230 796.000 27.510 800.000 ;
    END
  END input_pc[0]
  PIN input_pc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 524.030 796.000 524.310 800.000 ;
    END
  END input_pc[10]
  PIN input_pc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 573.710 796.000 573.990 800.000 ;
    END
  END input_pc[11]
  PIN input_pc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 623.390 796.000 623.670 800.000 ;
    END
  END input_pc[12]
  PIN input_pc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 673.070 796.000 673.350 800.000 ;
    END
  END input_pc[13]
  PIN input_pc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 722.750 796.000 723.030 800.000 ;
    END
  END input_pc[14]
  PIN input_pc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 772.430 796.000 772.710 800.000 ;
    END
  END input_pc[15]
  PIN input_pc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 76.910 796.000 77.190 800.000 ;
    END
  END input_pc[1]
  PIN input_pc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 126.590 796.000 126.870 800.000 ;
    END
  END input_pc[2]
  PIN input_pc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 176.270 796.000 176.550 800.000 ;
    END
  END input_pc[3]
  PIN input_pc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 225.950 796.000 226.230 800.000 ;
    END
  END input_pc[4]
  PIN input_pc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 275.630 796.000 275.910 800.000 ;
    END
  END input_pc[5]
  PIN input_pc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 325.310 796.000 325.590 800.000 ;
    END
  END input_pc[6]
  PIN input_pc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 374.990 796.000 375.270 800.000 ;
    END
  END input_pc[7]
  PIN input_pc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 424.670 796.000 424.950 800.000 ;
    END
  END input_pc[8]
  PIN input_pc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 474.350 796.000 474.630 800.000 ;
    END
  END input_pc[9]
  PIN output_ai[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END output_ai[0]
  PIN output_ai[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 4.000 ;
    END
  END output_ai[100]
  PIN output_ai[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END output_ai[101]
  PIN output_ai[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END output_ai[102]
  PIN output_ai[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END output_ai[103]
  PIN output_ai[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END output_ai[104]
  PIN output_ai[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 352.910 0.000 353.190 4.000 ;
    END
  END output_ai[105]
  PIN output_ai[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END output_ai[106]
  PIN output_ai[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END output_ai[107]
  PIN output_ai[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END output_ai[108]
  PIN output_ai[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END output_ai[109]
  PIN output_ai[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END output_ai[10]
  PIN output_ai[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END output_ai[110]
  PIN output_ai[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END output_ai[111]
  PIN output_ai[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END output_ai[112]
  PIN output_ai[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END output_ai[113]
  PIN output_ai[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 4.000 ;
    END
  END output_ai[114]
  PIN output_ai[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END output_ai[115]
  PIN output_ai[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END output_ai[116]
  PIN output_ai[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END output_ai[117]
  PIN output_ai[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END output_ai[118]
  PIN output_ai[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END output_ai[119]
  PIN output_ai[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END output_ai[11]
  PIN output_ai[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END output_ai[120]
  PIN output_ai[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END output_ai[121]
  PIN output_ai[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END output_ai[122]
  PIN output_ai[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END output_ai[123]
  PIN output_ai[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 4.000 ;
    END
  END output_ai[124]
  PIN output_ai[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END output_ai[125]
  PIN output_ai[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END output_ai[126]
  PIN output_ai[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END output_ai[127]
  PIN output_ai[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END output_ai[128]
  PIN output_ai[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END output_ai[129]
  PIN output_ai[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END output_ai[12]
  PIN output_ai[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END output_ai[130]
  PIN output_ai[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 436.630 0.000 436.910 4.000 ;
    END
  END output_ai[131]
  PIN output_ai[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 439.850 0.000 440.130 4.000 ;
    END
  END output_ai[132]
  PIN output_ai[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END output_ai[133]
  PIN output_ai[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END output_ai[134]
  PIN output_ai[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END output_ai[135]
  PIN output_ai[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END output_ai[136]
  PIN output_ai[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 455.950 0.000 456.230 4.000 ;
    END
  END output_ai[137]
  PIN output_ai[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 459.170 0.000 459.450 4.000 ;
    END
  END output_ai[138]
  PIN output_ai[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END output_ai[139]
  PIN output_ai[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END output_ai[13]
  PIN output_ai[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END output_ai[140]
  PIN output_ai[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 468.830 0.000 469.110 4.000 ;
    END
  END output_ai[141]
  PIN output_ai[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END output_ai[142]
  PIN output_ai[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END output_ai[143]
  PIN output_ai[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END output_ai[144]
  PIN output_ai[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END output_ai[145]
  PIN output_ai[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END output_ai[146]
  PIN output_ai[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END output_ai[147]
  PIN output_ai[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END output_ai[148]
  PIN output_ai[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END output_ai[149]
  PIN output_ai[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END output_ai[14]
  PIN output_ai[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END output_ai[150]
  PIN output_ai[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END output_ai[151]
  PIN output_ai[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END output_ai[152]
  PIN output_ai[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END output_ai[153]
  PIN output_ai[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END output_ai[154]
  PIN output_ai[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END output_ai[155]
  PIN output_ai[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END output_ai[156]
  PIN output_ai[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END output_ai[157]
  PIN output_ai[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END output_ai[158]
  PIN output_ai[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END output_ai[159]
  PIN output_ai[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END output_ai[15]
  PIN output_ai[160]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END output_ai[160]
  PIN output_ai[161]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END output_ai[161]
  PIN output_ai[162]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END output_ai[162]
  PIN output_ai[163]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END output_ai[163]
  PIN output_ai[164]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END output_ai[164]
  PIN output_ai[165]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END output_ai[165]
  PIN output_ai[166]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END output_ai[166]
  PIN output_ai[167]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END output_ai[167]
  PIN output_ai[168]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END output_ai[168]
  PIN output_ai[169]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END output_ai[169]
  PIN output_ai[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END output_ai[16]
  PIN output_ai[170]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END output_ai[170]
  PIN output_ai[171]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 565.430 0.000 565.710 4.000 ;
    END
  END output_ai[171]
  PIN output_ai[172]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END output_ai[172]
  PIN output_ai[173]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END output_ai[173]
  PIN output_ai[174]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END output_ai[174]
  PIN output_ai[175]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END output_ai[175]
  PIN output_ai[176]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END output_ai[176]
  PIN output_ai[177]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 584.750 0.000 585.030 4.000 ;
    END
  END output_ai[177]
  PIN output_ai[178]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END output_ai[178]
  PIN output_ai[179]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 591.190 0.000 591.470 4.000 ;
    END
  END output_ai[179]
  PIN output_ai[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END output_ai[17]
  PIN output_ai[180]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 594.410 0.000 594.690 4.000 ;
    END
  END output_ai[180]
  PIN output_ai[181]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END output_ai[181]
  PIN output_ai[182]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END output_ai[182]
  PIN output_ai[183]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END output_ai[183]
  PIN output_ai[184]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END output_ai[184]
  PIN output_ai[185]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END output_ai[185]
  PIN output_ai[186]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 4.000 ;
    END
  END output_ai[186]
  PIN output_ai[187]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END output_ai[187]
  PIN output_ai[188]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END output_ai[188]
  PIN output_ai[189]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END output_ai[189]
  PIN output_ai[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END output_ai[18]
  PIN output_ai[190]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END output_ai[190]
  PIN output_ai[191]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END output_ai[191]
  PIN output_ai[192]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END output_ai[192]
  PIN output_ai[193]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END output_ai[193]
  PIN output_ai[194]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END output_ai[194]
  PIN output_ai[195]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END output_ai[195]
  PIN output_ai[196]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END output_ai[196]
  PIN output_ai[197]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END output_ai[197]
  PIN output_ai[198]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END output_ai[198]
  PIN output_ai[199]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END output_ai[199]
  PIN output_ai[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END output_ai[19]
  PIN output_ai[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END output_ai[1]
  PIN output_ai[200]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 658.810 0.000 659.090 4.000 ;
    END
  END output_ai[200]
  PIN output_ai[201]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 662.030 0.000 662.310 4.000 ;
    END
  END output_ai[201]
  PIN output_ai[202]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END output_ai[202]
  PIN output_ai[203]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 4.000 ;
    END
  END output_ai[203]
  PIN output_ai[204]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END output_ai[204]
  PIN output_ai[205]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END output_ai[205]
  PIN output_ai[206]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 678.130 0.000 678.410 4.000 ;
    END
  END output_ai[206]
  PIN output_ai[207]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END output_ai[207]
  PIN output_ai[208]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END output_ai[208]
  PIN output_ai[209]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END output_ai[209]
  PIN output_ai[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END output_ai[20]
  PIN output_ai[210]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END output_ai[210]
  PIN output_ai[211]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END output_ai[211]
  PIN output_ai[212]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END output_ai[212]
  PIN output_ai[213]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END output_ai[213]
  PIN output_ai[214]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 703.890 0.000 704.170 4.000 ;
    END
  END output_ai[214]
  PIN output_ai[215]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 4.000 ;
    END
  END output_ai[215]
  PIN output_ai[216]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END output_ai[216]
  PIN output_ai[217]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END output_ai[217]
  PIN output_ai[218]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END output_ai[218]
  PIN output_ai[219]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END output_ai[219]
  PIN output_ai[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END output_ai[21]
  PIN output_ai[220]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 4.000 ;
    END
  END output_ai[220]
  PIN output_ai[221]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END output_ai[221]
  PIN output_ai[222]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END output_ai[222]
  PIN output_ai[223]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END output_ai[223]
  PIN output_ai[224]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END output_ai[224]
  PIN output_ai[225]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 739.310 0.000 739.590 4.000 ;
    END
  END output_ai[225]
  PIN output_ai[226]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END output_ai[226]
  PIN output_ai[227]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 745.750 0.000 746.030 4.000 ;
    END
  END output_ai[227]
  PIN output_ai[228]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 748.970 0.000 749.250 4.000 ;
    END
  END output_ai[228]
  PIN output_ai[229]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END output_ai[229]
  PIN output_ai[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END output_ai[22]
  PIN output_ai[230]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END output_ai[230]
  PIN output_ai[231]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END output_ai[231]
  PIN output_ai[232]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 761.850 0.000 762.130 4.000 ;
    END
  END output_ai[232]
  PIN output_ai[233]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 765.070 0.000 765.350 4.000 ;
    END
  END output_ai[233]
  PIN output_ai[234]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END output_ai[234]
  PIN output_ai[235]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END output_ai[235]
  PIN output_ai[236]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END output_ai[236]
  PIN output_ai[237]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END output_ai[237]
  PIN output_ai[238]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END output_ai[238]
  PIN output_ai[239]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END output_ai[239]
  PIN output_ai[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END output_ai[23]
  PIN output_ai[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END output_ai[24]
  PIN output_ai[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END output_ai[25]
  PIN output_ai[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END output_ai[26]
  PIN output_ai[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END output_ai[27]
  PIN output_ai[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END output_ai[28]
  PIN output_ai[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END output_ai[29]
  PIN output_ai[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END output_ai[2]
  PIN output_ai[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END output_ai[30]
  PIN output_ai[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END output_ai[31]
  PIN output_ai[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END output_ai[32]
  PIN output_ai[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END output_ai[33]
  PIN output_ai[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END output_ai[34]
  PIN output_ai[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END output_ai[35]
  PIN output_ai[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END output_ai[36]
  PIN output_ai[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END output_ai[37]
  PIN output_ai[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END output_ai[38]
  PIN output_ai[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END output_ai[39]
  PIN output_ai[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END output_ai[3]
  PIN output_ai[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END output_ai[40]
  PIN output_ai[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 146.830 0.000 147.110 4.000 ;
    END
  END output_ai[41]
  PIN output_ai[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END output_ai[42]
  PIN output_ai[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END output_ai[43]
  PIN output_ai[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END output_ai[44]
  PIN output_ai[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 159.710 0.000 159.990 4.000 ;
    END
  END output_ai[45]
  PIN output_ai[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END output_ai[46]
  PIN output_ai[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END output_ai[47]
  PIN output_ai[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END output_ai[48]
  PIN output_ai[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END output_ai[49]
  PIN output_ai[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END output_ai[4]
  PIN output_ai[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END output_ai[50]
  PIN output_ai[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END output_ai[51]
  PIN output_ai[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END output_ai[52]
  PIN output_ai[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END output_ai[53]
  PIN output_ai[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END output_ai[54]
  PIN output_ai[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END output_ai[55]
  PIN output_ai[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END output_ai[56]
  PIN output_ai[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END output_ai[57]
  PIN output_ai[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END output_ai[58]
  PIN output_ai[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 204.790 0.000 205.070 4.000 ;
    END
  END output_ai[59]
  PIN output_ai[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END output_ai[5]
  PIN output_ai[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END output_ai[60]
  PIN output_ai[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 211.230 0.000 211.510 4.000 ;
    END
  END output_ai[61]
  PIN output_ai[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END output_ai[62]
  PIN output_ai[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END output_ai[63]
  PIN output_ai[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END output_ai[64]
  PIN output_ai[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 224.110 0.000 224.390 4.000 ;
    END
  END output_ai[65]
  PIN output_ai[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 227.330 0.000 227.610 4.000 ;
    END
  END output_ai[66]
  PIN output_ai[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END output_ai[67]
  PIN output_ai[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END output_ai[68]
  PIN output_ai[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END output_ai[69]
  PIN output_ai[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END output_ai[6]
  PIN output_ai[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END output_ai[70]
  PIN output_ai[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END output_ai[71]
  PIN output_ai[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END output_ai[72]
  PIN output_ai[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END output_ai[73]
  PIN output_ai[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END output_ai[74]
  PIN output_ai[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END output_ai[75]
  PIN output_ai[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END output_ai[76]
  PIN output_ai[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END output_ai[77]
  PIN output_ai[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 265.970 0.000 266.250 4.000 ;
    END
  END output_ai[78]
  PIN output_ai[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 4.000 ;
    END
  END output_ai[79]
  PIN output_ai[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END output_ai[7]
  PIN output_ai[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END output_ai[80]
  PIN output_ai[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END output_ai[81]
  PIN output_ai[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END output_ai[82]
  PIN output_ai[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END output_ai[83]
  PIN output_ai[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 285.290 0.000 285.570 4.000 ;
    END
  END output_ai[84]
  PIN output_ai[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 288.510 0.000 288.790 4.000 ;
    END
  END output_ai[85]
  PIN output_ai[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END output_ai[86]
  PIN output_ai[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END output_ai[87]
  PIN output_ai[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END output_ai[88]
  PIN output_ai[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END output_ai[89]
  PIN output_ai[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END output_ai[8]
  PIN output_ai[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END output_ai[90]
  PIN output_ai[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END output_ai[91]
  PIN output_ai[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END output_ai[92]
  PIN output_ai[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END output_ai[93]
  PIN output_ai[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END output_ai[94]
  PIN output_ai[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END output_ai[95]
  PIN output_ai[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END output_ai[96]
  PIN output_ai[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END output_ai[97]
  PIN output_ai[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END output_ai[98]
  PIN output_ai[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END output_ai[99]
  PIN output_ai[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END output_ai[9]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END reset
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 788.885 ;
      LAYER met1 ;
        RECT 5.520 9.900 794.420 789.040 ;
      LAYER met2 ;
        RECT 7.450 795.720 26.950 796.690 ;
        RECT 27.790 795.720 76.630 796.690 ;
        RECT 77.470 795.720 126.310 796.690 ;
        RECT 127.150 795.720 175.990 796.690 ;
        RECT 176.830 795.720 225.670 796.690 ;
        RECT 226.510 795.720 275.350 796.690 ;
        RECT 276.190 795.720 325.030 796.690 ;
        RECT 325.870 795.720 374.710 796.690 ;
        RECT 375.550 795.720 424.390 796.690 ;
        RECT 425.230 795.720 474.070 796.690 ;
        RECT 474.910 795.720 523.750 796.690 ;
        RECT 524.590 795.720 573.430 796.690 ;
        RECT 574.270 795.720 623.110 796.690 ;
        RECT 623.950 795.720 672.790 796.690 ;
        RECT 673.630 795.720 722.470 796.690 ;
        RECT 723.310 795.720 772.150 796.690 ;
        RECT 772.990 795.720 793.910 796.690 ;
        RECT 7.450 4.280 793.910 795.720 ;
        RECT 7.450 3.670 14.530 4.280 ;
        RECT 15.370 3.670 17.750 4.280 ;
        RECT 18.590 3.670 20.970 4.280 ;
        RECT 21.810 3.670 24.190 4.280 ;
        RECT 25.030 3.670 27.410 4.280 ;
        RECT 28.250 3.670 30.630 4.280 ;
        RECT 31.470 3.670 33.850 4.280 ;
        RECT 34.690 3.670 37.070 4.280 ;
        RECT 37.910 3.670 40.290 4.280 ;
        RECT 41.130 3.670 43.510 4.280 ;
        RECT 44.350 3.670 46.730 4.280 ;
        RECT 47.570 3.670 49.950 4.280 ;
        RECT 50.790 3.670 53.170 4.280 ;
        RECT 54.010 3.670 56.390 4.280 ;
        RECT 57.230 3.670 59.610 4.280 ;
        RECT 60.450 3.670 62.830 4.280 ;
        RECT 63.670 3.670 66.050 4.280 ;
        RECT 66.890 3.670 69.270 4.280 ;
        RECT 70.110 3.670 72.490 4.280 ;
        RECT 73.330 3.670 75.710 4.280 ;
        RECT 76.550 3.670 78.930 4.280 ;
        RECT 79.770 3.670 82.150 4.280 ;
        RECT 82.990 3.670 85.370 4.280 ;
        RECT 86.210 3.670 88.590 4.280 ;
        RECT 89.430 3.670 91.810 4.280 ;
        RECT 92.650 3.670 95.030 4.280 ;
        RECT 95.870 3.670 98.250 4.280 ;
        RECT 99.090 3.670 101.470 4.280 ;
        RECT 102.310 3.670 104.690 4.280 ;
        RECT 105.530 3.670 107.910 4.280 ;
        RECT 108.750 3.670 111.130 4.280 ;
        RECT 111.970 3.670 114.350 4.280 ;
        RECT 115.190 3.670 117.570 4.280 ;
        RECT 118.410 3.670 120.790 4.280 ;
        RECT 121.630 3.670 124.010 4.280 ;
        RECT 124.850 3.670 127.230 4.280 ;
        RECT 128.070 3.670 130.450 4.280 ;
        RECT 131.290 3.670 133.670 4.280 ;
        RECT 134.510 3.670 136.890 4.280 ;
        RECT 137.730 3.670 140.110 4.280 ;
        RECT 140.950 3.670 143.330 4.280 ;
        RECT 144.170 3.670 146.550 4.280 ;
        RECT 147.390 3.670 149.770 4.280 ;
        RECT 150.610 3.670 152.990 4.280 ;
        RECT 153.830 3.670 156.210 4.280 ;
        RECT 157.050 3.670 159.430 4.280 ;
        RECT 160.270 3.670 162.650 4.280 ;
        RECT 163.490 3.670 165.870 4.280 ;
        RECT 166.710 3.670 169.090 4.280 ;
        RECT 169.930 3.670 172.310 4.280 ;
        RECT 173.150 3.670 175.530 4.280 ;
        RECT 176.370 3.670 178.750 4.280 ;
        RECT 179.590 3.670 181.970 4.280 ;
        RECT 182.810 3.670 185.190 4.280 ;
        RECT 186.030 3.670 188.410 4.280 ;
        RECT 189.250 3.670 191.630 4.280 ;
        RECT 192.470 3.670 194.850 4.280 ;
        RECT 195.690 3.670 198.070 4.280 ;
        RECT 198.910 3.670 201.290 4.280 ;
        RECT 202.130 3.670 204.510 4.280 ;
        RECT 205.350 3.670 207.730 4.280 ;
        RECT 208.570 3.670 210.950 4.280 ;
        RECT 211.790 3.670 214.170 4.280 ;
        RECT 215.010 3.670 217.390 4.280 ;
        RECT 218.230 3.670 220.610 4.280 ;
        RECT 221.450 3.670 223.830 4.280 ;
        RECT 224.670 3.670 227.050 4.280 ;
        RECT 227.890 3.670 230.270 4.280 ;
        RECT 231.110 3.670 233.490 4.280 ;
        RECT 234.330 3.670 236.710 4.280 ;
        RECT 237.550 3.670 239.930 4.280 ;
        RECT 240.770 3.670 243.150 4.280 ;
        RECT 243.990 3.670 246.370 4.280 ;
        RECT 247.210 3.670 249.590 4.280 ;
        RECT 250.430 3.670 252.810 4.280 ;
        RECT 253.650 3.670 256.030 4.280 ;
        RECT 256.870 3.670 259.250 4.280 ;
        RECT 260.090 3.670 262.470 4.280 ;
        RECT 263.310 3.670 265.690 4.280 ;
        RECT 266.530 3.670 268.910 4.280 ;
        RECT 269.750 3.670 272.130 4.280 ;
        RECT 272.970 3.670 275.350 4.280 ;
        RECT 276.190 3.670 278.570 4.280 ;
        RECT 279.410 3.670 281.790 4.280 ;
        RECT 282.630 3.670 285.010 4.280 ;
        RECT 285.850 3.670 288.230 4.280 ;
        RECT 289.070 3.670 291.450 4.280 ;
        RECT 292.290 3.670 294.670 4.280 ;
        RECT 295.510 3.670 297.890 4.280 ;
        RECT 298.730 3.670 301.110 4.280 ;
        RECT 301.950 3.670 304.330 4.280 ;
        RECT 305.170 3.670 307.550 4.280 ;
        RECT 308.390 3.670 310.770 4.280 ;
        RECT 311.610 3.670 313.990 4.280 ;
        RECT 314.830 3.670 317.210 4.280 ;
        RECT 318.050 3.670 320.430 4.280 ;
        RECT 321.270 3.670 323.650 4.280 ;
        RECT 324.490 3.670 326.870 4.280 ;
        RECT 327.710 3.670 330.090 4.280 ;
        RECT 330.930 3.670 333.310 4.280 ;
        RECT 334.150 3.670 336.530 4.280 ;
        RECT 337.370 3.670 339.750 4.280 ;
        RECT 340.590 3.670 342.970 4.280 ;
        RECT 343.810 3.670 346.190 4.280 ;
        RECT 347.030 3.670 349.410 4.280 ;
        RECT 350.250 3.670 352.630 4.280 ;
        RECT 353.470 3.670 355.850 4.280 ;
        RECT 356.690 3.670 359.070 4.280 ;
        RECT 359.910 3.670 362.290 4.280 ;
        RECT 363.130 3.670 365.510 4.280 ;
        RECT 366.350 3.670 368.730 4.280 ;
        RECT 369.570 3.670 371.950 4.280 ;
        RECT 372.790 3.670 375.170 4.280 ;
        RECT 376.010 3.670 378.390 4.280 ;
        RECT 379.230 3.670 381.610 4.280 ;
        RECT 382.450 3.670 384.830 4.280 ;
        RECT 385.670 3.670 388.050 4.280 ;
        RECT 388.890 3.670 391.270 4.280 ;
        RECT 392.110 3.670 394.490 4.280 ;
        RECT 395.330 3.670 397.710 4.280 ;
        RECT 398.550 3.670 400.930 4.280 ;
        RECT 401.770 3.670 404.150 4.280 ;
        RECT 404.990 3.670 407.370 4.280 ;
        RECT 408.210 3.670 410.590 4.280 ;
        RECT 411.430 3.670 413.810 4.280 ;
        RECT 414.650 3.670 417.030 4.280 ;
        RECT 417.870 3.670 420.250 4.280 ;
        RECT 421.090 3.670 423.470 4.280 ;
        RECT 424.310 3.670 426.690 4.280 ;
        RECT 427.530 3.670 429.910 4.280 ;
        RECT 430.750 3.670 433.130 4.280 ;
        RECT 433.970 3.670 436.350 4.280 ;
        RECT 437.190 3.670 439.570 4.280 ;
        RECT 440.410 3.670 442.790 4.280 ;
        RECT 443.630 3.670 446.010 4.280 ;
        RECT 446.850 3.670 449.230 4.280 ;
        RECT 450.070 3.670 452.450 4.280 ;
        RECT 453.290 3.670 455.670 4.280 ;
        RECT 456.510 3.670 458.890 4.280 ;
        RECT 459.730 3.670 462.110 4.280 ;
        RECT 462.950 3.670 465.330 4.280 ;
        RECT 466.170 3.670 468.550 4.280 ;
        RECT 469.390 3.670 471.770 4.280 ;
        RECT 472.610 3.670 474.990 4.280 ;
        RECT 475.830 3.670 478.210 4.280 ;
        RECT 479.050 3.670 481.430 4.280 ;
        RECT 482.270 3.670 484.650 4.280 ;
        RECT 485.490 3.670 487.870 4.280 ;
        RECT 488.710 3.670 491.090 4.280 ;
        RECT 491.930 3.670 494.310 4.280 ;
        RECT 495.150 3.670 497.530 4.280 ;
        RECT 498.370 3.670 500.750 4.280 ;
        RECT 501.590 3.670 503.970 4.280 ;
        RECT 504.810 3.670 507.190 4.280 ;
        RECT 508.030 3.670 510.410 4.280 ;
        RECT 511.250 3.670 513.630 4.280 ;
        RECT 514.470 3.670 516.850 4.280 ;
        RECT 517.690 3.670 520.070 4.280 ;
        RECT 520.910 3.670 523.290 4.280 ;
        RECT 524.130 3.670 526.510 4.280 ;
        RECT 527.350 3.670 529.730 4.280 ;
        RECT 530.570 3.670 532.950 4.280 ;
        RECT 533.790 3.670 536.170 4.280 ;
        RECT 537.010 3.670 539.390 4.280 ;
        RECT 540.230 3.670 542.610 4.280 ;
        RECT 543.450 3.670 545.830 4.280 ;
        RECT 546.670 3.670 549.050 4.280 ;
        RECT 549.890 3.670 552.270 4.280 ;
        RECT 553.110 3.670 555.490 4.280 ;
        RECT 556.330 3.670 558.710 4.280 ;
        RECT 559.550 3.670 561.930 4.280 ;
        RECT 562.770 3.670 565.150 4.280 ;
        RECT 565.990 3.670 568.370 4.280 ;
        RECT 569.210 3.670 571.590 4.280 ;
        RECT 572.430 3.670 574.810 4.280 ;
        RECT 575.650 3.670 578.030 4.280 ;
        RECT 578.870 3.670 581.250 4.280 ;
        RECT 582.090 3.670 584.470 4.280 ;
        RECT 585.310 3.670 587.690 4.280 ;
        RECT 588.530 3.670 590.910 4.280 ;
        RECT 591.750 3.670 594.130 4.280 ;
        RECT 594.970 3.670 597.350 4.280 ;
        RECT 598.190 3.670 600.570 4.280 ;
        RECT 601.410 3.670 603.790 4.280 ;
        RECT 604.630 3.670 607.010 4.280 ;
        RECT 607.850 3.670 610.230 4.280 ;
        RECT 611.070 3.670 613.450 4.280 ;
        RECT 614.290 3.670 616.670 4.280 ;
        RECT 617.510 3.670 619.890 4.280 ;
        RECT 620.730 3.670 623.110 4.280 ;
        RECT 623.950 3.670 626.330 4.280 ;
        RECT 627.170 3.670 629.550 4.280 ;
        RECT 630.390 3.670 632.770 4.280 ;
        RECT 633.610 3.670 635.990 4.280 ;
        RECT 636.830 3.670 639.210 4.280 ;
        RECT 640.050 3.670 642.430 4.280 ;
        RECT 643.270 3.670 645.650 4.280 ;
        RECT 646.490 3.670 648.870 4.280 ;
        RECT 649.710 3.670 652.090 4.280 ;
        RECT 652.930 3.670 655.310 4.280 ;
        RECT 656.150 3.670 658.530 4.280 ;
        RECT 659.370 3.670 661.750 4.280 ;
        RECT 662.590 3.670 664.970 4.280 ;
        RECT 665.810 3.670 668.190 4.280 ;
        RECT 669.030 3.670 671.410 4.280 ;
        RECT 672.250 3.670 674.630 4.280 ;
        RECT 675.470 3.670 677.850 4.280 ;
        RECT 678.690 3.670 681.070 4.280 ;
        RECT 681.910 3.670 684.290 4.280 ;
        RECT 685.130 3.670 687.510 4.280 ;
        RECT 688.350 3.670 690.730 4.280 ;
        RECT 691.570 3.670 693.950 4.280 ;
        RECT 694.790 3.670 697.170 4.280 ;
        RECT 698.010 3.670 700.390 4.280 ;
        RECT 701.230 3.670 703.610 4.280 ;
        RECT 704.450 3.670 706.830 4.280 ;
        RECT 707.670 3.670 710.050 4.280 ;
        RECT 710.890 3.670 713.270 4.280 ;
        RECT 714.110 3.670 716.490 4.280 ;
        RECT 717.330 3.670 719.710 4.280 ;
        RECT 720.550 3.670 722.930 4.280 ;
        RECT 723.770 3.670 726.150 4.280 ;
        RECT 726.990 3.670 729.370 4.280 ;
        RECT 730.210 3.670 732.590 4.280 ;
        RECT 733.430 3.670 735.810 4.280 ;
        RECT 736.650 3.670 739.030 4.280 ;
        RECT 739.870 3.670 742.250 4.280 ;
        RECT 743.090 3.670 745.470 4.280 ;
        RECT 746.310 3.670 748.690 4.280 ;
        RECT 749.530 3.670 751.910 4.280 ;
        RECT 752.750 3.670 755.130 4.280 ;
        RECT 755.970 3.670 758.350 4.280 ;
        RECT 759.190 3.670 761.570 4.280 ;
        RECT 762.410 3.670 764.790 4.280 ;
        RECT 765.630 3.670 768.010 4.280 ;
        RECT 768.850 3.670 771.230 4.280 ;
        RECT 772.070 3.670 774.450 4.280 ;
        RECT 775.290 3.670 777.670 4.280 ;
        RECT 778.510 3.670 780.890 4.280 ;
        RECT 781.730 3.670 784.110 4.280 ;
        RECT 784.950 3.670 793.910 4.280 ;
      LAYER met3 ;
        RECT 4.000 399.520 796.000 788.965 ;
        RECT 4.400 398.120 795.600 399.520 ;
        RECT 4.000 10.715 796.000 398.120 ;
  END
END shifter
END LIBRARY

