VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO lowpass
  CLASS BLOCK ;
  FOREIGN lowpass ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.540 10.640 333.140 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 485.140 10.640 486.740 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.740 10.640 640.340 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 792.340 10.640 793.940 789.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 796.000 398.520 800.000 399.120 ;
    END
  END clk
  PIN input_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 14.810 796.000 15.090 800.000 ;
    END
  END input_data[0]
  PIN input_data[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 336.810 796.000 337.090 800.000 ;
    END
  END input_data[100]
  PIN input_data[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 340.030 796.000 340.310 800.000 ;
    END
  END input_data[101]
  PIN input_data[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 343.250 796.000 343.530 800.000 ;
    END
  END input_data[102]
  PIN input_data[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 346.470 796.000 346.750 800.000 ;
    END
  END input_data[103]
  PIN input_data[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.690 796.000 349.970 800.000 ;
    END
  END input_data[104]
  PIN input_data[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 352.910 796.000 353.190 800.000 ;
    END
  END input_data[105]
  PIN input_data[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 356.130 796.000 356.410 800.000 ;
    END
  END input_data[106]
  PIN input_data[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 359.350 796.000 359.630 800.000 ;
    END
  END input_data[107]
  PIN input_data[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 362.570 796.000 362.850 800.000 ;
    END
  END input_data[108]
  PIN input_data[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 365.790 796.000 366.070 800.000 ;
    END
  END input_data[109]
  PIN input_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 47.010 796.000 47.290 800.000 ;
    END
  END input_data[10]
  PIN input_data[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 369.010 796.000 369.290 800.000 ;
    END
  END input_data[110]
  PIN input_data[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 372.230 796.000 372.510 800.000 ;
    END
  END input_data[111]
  PIN input_data[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 375.450 796.000 375.730 800.000 ;
    END
  END input_data[112]
  PIN input_data[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 378.670 796.000 378.950 800.000 ;
    END
  END input_data[113]
  PIN input_data[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 381.890 796.000 382.170 800.000 ;
    END
  END input_data[114]
  PIN input_data[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 385.110 796.000 385.390 800.000 ;
    END
  END input_data[115]
  PIN input_data[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 388.330 796.000 388.610 800.000 ;
    END
  END input_data[116]
  PIN input_data[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 391.550 796.000 391.830 800.000 ;
    END
  END input_data[117]
  PIN input_data[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 394.770 796.000 395.050 800.000 ;
    END
  END input_data[118]
  PIN input_data[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 397.990 796.000 398.270 800.000 ;
    END
  END input_data[119]
  PIN input_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 50.230 796.000 50.510 800.000 ;
    END
  END input_data[11]
  PIN input_data[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 401.210 796.000 401.490 800.000 ;
    END
  END input_data[120]
  PIN input_data[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 404.430 796.000 404.710 800.000 ;
    END
  END input_data[121]
  PIN input_data[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 407.650 796.000 407.930 800.000 ;
    END
  END input_data[122]
  PIN input_data[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 410.870 796.000 411.150 800.000 ;
    END
  END input_data[123]
  PIN input_data[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 414.090 796.000 414.370 800.000 ;
    END
  END input_data[124]
  PIN input_data[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 417.310 796.000 417.590 800.000 ;
    END
  END input_data[125]
  PIN input_data[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 420.530 796.000 420.810 800.000 ;
    END
  END input_data[126]
  PIN input_data[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 423.750 796.000 424.030 800.000 ;
    END
  END input_data[127]
  PIN input_data[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 426.970 796.000 427.250 800.000 ;
    END
  END input_data[128]
  PIN input_data[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 430.190 796.000 430.470 800.000 ;
    END
  END input_data[129]
  PIN input_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.450 796.000 53.730 800.000 ;
    END
  END input_data[12]
  PIN input_data[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 433.410 796.000 433.690 800.000 ;
    END
  END input_data[130]
  PIN input_data[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 436.630 796.000 436.910 800.000 ;
    END
  END input_data[131]
  PIN input_data[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 439.850 796.000 440.130 800.000 ;
    END
  END input_data[132]
  PIN input_data[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 443.070 796.000 443.350 800.000 ;
    END
  END input_data[133]
  PIN input_data[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 446.290 796.000 446.570 800.000 ;
    END
  END input_data[134]
  PIN input_data[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 449.510 796.000 449.790 800.000 ;
    END
  END input_data[135]
  PIN input_data[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 452.730 796.000 453.010 800.000 ;
    END
  END input_data[136]
  PIN input_data[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 455.950 796.000 456.230 800.000 ;
    END
  END input_data[137]
  PIN input_data[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 459.170 796.000 459.450 800.000 ;
    END
  END input_data[138]
  PIN input_data[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 462.390 796.000 462.670 800.000 ;
    END
  END input_data[139]
  PIN input_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.670 796.000 56.950 800.000 ;
    END
  END input_data[13]
  PIN input_data[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 465.610 796.000 465.890 800.000 ;
    END
  END input_data[140]
  PIN input_data[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 468.830 796.000 469.110 800.000 ;
    END
  END input_data[141]
  PIN input_data[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 472.050 796.000 472.330 800.000 ;
    END
  END input_data[142]
  PIN input_data[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 475.270 796.000 475.550 800.000 ;
    END
  END input_data[143]
  PIN input_data[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 478.490 796.000 478.770 800.000 ;
    END
  END input_data[144]
  PIN input_data[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 481.710 796.000 481.990 800.000 ;
    END
  END input_data[145]
  PIN input_data[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 484.930 796.000 485.210 800.000 ;
    END
  END input_data[146]
  PIN input_data[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 488.150 796.000 488.430 800.000 ;
    END
  END input_data[147]
  PIN input_data[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 491.370 796.000 491.650 800.000 ;
    END
  END input_data[148]
  PIN input_data[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 494.590 796.000 494.870 800.000 ;
    END
  END input_data[149]
  PIN input_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.890 796.000 60.170 800.000 ;
    END
  END input_data[14]
  PIN input_data[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 497.810 796.000 498.090 800.000 ;
    END
  END input_data[150]
  PIN input_data[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 501.030 796.000 501.310 800.000 ;
    END
  END input_data[151]
  PIN input_data[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 504.250 796.000 504.530 800.000 ;
    END
  END input_data[152]
  PIN input_data[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 507.470 796.000 507.750 800.000 ;
    END
  END input_data[153]
  PIN input_data[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 510.690 796.000 510.970 800.000 ;
    END
  END input_data[154]
  PIN input_data[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 513.910 796.000 514.190 800.000 ;
    END
  END input_data[155]
  PIN input_data[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 517.130 796.000 517.410 800.000 ;
    END
  END input_data[156]
  PIN input_data[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 520.350 796.000 520.630 800.000 ;
    END
  END input_data[157]
  PIN input_data[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 523.570 796.000 523.850 800.000 ;
    END
  END input_data[158]
  PIN input_data[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 526.790 796.000 527.070 800.000 ;
    END
  END input_data[159]
  PIN input_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 796.000 63.390 800.000 ;
    END
  END input_data[15]
  PIN input_data[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 530.010 796.000 530.290 800.000 ;
    END
  END input_data[160]
  PIN input_data[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 533.230 796.000 533.510 800.000 ;
    END
  END input_data[161]
  PIN input_data[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 536.450 796.000 536.730 800.000 ;
    END
  END input_data[162]
  PIN input_data[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 539.670 796.000 539.950 800.000 ;
    END
  END input_data[163]
  PIN input_data[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 542.890 796.000 543.170 800.000 ;
    END
  END input_data[164]
  PIN input_data[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 546.110 796.000 546.390 800.000 ;
    END
  END input_data[165]
  PIN input_data[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 549.330 796.000 549.610 800.000 ;
    END
  END input_data[166]
  PIN input_data[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 552.550 796.000 552.830 800.000 ;
    END
  END input_data[167]
  PIN input_data[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 555.770 796.000 556.050 800.000 ;
    END
  END input_data[168]
  PIN input_data[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 558.990 796.000 559.270 800.000 ;
    END
  END input_data[169]
  PIN input_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 66.330 796.000 66.610 800.000 ;
    END
  END input_data[16]
  PIN input_data[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 562.210 796.000 562.490 800.000 ;
    END
  END input_data[170]
  PIN input_data[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 565.430 796.000 565.710 800.000 ;
    END
  END input_data[171]
  PIN input_data[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 568.650 796.000 568.930 800.000 ;
    END
  END input_data[172]
  PIN input_data[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 571.870 796.000 572.150 800.000 ;
    END
  END input_data[173]
  PIN input_data[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 575.090 796.000 575.370 800.000 ;
    END
  END input_data[174]
  PIN input_data[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 796.000 578.590 800.000 ;
    END
  END input_data[175]
  PIN input_data[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 581.530 796.000 581.810 800.000 ;
    END
  END input_data[176]
  PIN input_data[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 584.750 796.000 585.030 800.000 ;
    END
  END input_data[177]
  PIN input_data[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 587.970 796.000 588.250 800.000 ;
    END
  END input_data[178]
  PIN input_data[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 591.190 796.000 591.470 800.000 ;
    END
  END input_data[179]
  PIN input_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 69.550 796.000 69.830 800.000 ;
    END
  END input_data[17]
  PIN input_data[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 594.410 796.000 594.690 800.000 ;
    END
  END input_data[180]
  PIN input_data[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 597.630 796.000 597.910 800.000 ;
    END
  END input_data[181]
  PIN input_data[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 600.850 796.000 601.130 800.000 ;
    END
  END input_data[182]
  PIN input_data[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 604.070 796.000 604.350 800.000 ;
    END
  END input_data[183]
  PIN input_data[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 607.290 796.000 607.570 800.000 ;
    END
  END input_data[184]
  PIN input_data[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 610.510 796.000 610.790 800.000 ;
    END
  END input_data[185]
  PIN input_data[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 613.730 796.000 614.010 800.000 ;
    END
  END input_data[186]
  PIN input_data[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 616.950 796.000 617.230 800.000 ;
    END
  END input_data[187]
  PIN input_data[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 620.170 796.000 620.450 800.000 ;
    END
  END input_data[188]
  PIN input_data[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 623.390 796.000 623.670 800.000 ;
    END
  END input_data[189]
  PIN input_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 72.770 796.000 73.050 800.000 ;
    END
  END input_data[18]
  PIN input_data[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 626.610 796.000 626.890 800.000 ;
    END
  END input_data[190]
  PIN input_data[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 796.000 630.110 800.000 ;
    END
  END input_data[191]
  PIN input_data[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 633.050 796.000 633.330 800.000 ;
    END
  END input_data[192]
  PIN input_data[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 636.270 796.000 636.550 800.000 ;
    END
  END input_data[193]
  PIN input_data[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 639.490 796.000 639.770 800.000 ;
    END
  END input_data[194]
  PIN input_data[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 642.710 796.000 642.990 800.000 ;
    END
  END input_data[195]
  PIN input_data[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 645.930 796.000 646.210 800.000 ;
    END
  END input_data[196]
  PIN input_data[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 649.150 796.000 649.430 800.000 ;
    END
  END input_data[197]
  PIN input_data[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 652.370 796.000 652.650 800.000 ;
    END
  END input_data[198]
  PIN input_data[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 655.590 796.000 655.870 800.000 ;
    END
  END input_data[199]
  PIN input_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.990 796.000 76.270 800.000 ;
    END
  END input_data[19]
  PIN input_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 18.030 796.000 18.310 800.000 ;
    END
  END input_data[1]
  PIN input_data[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 658.810 796.000 659.090 800.000 ;
    END
  END input_data[200]
  PIN input_data[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 662.030 796.000 662.310 800.000 ;
    END
  END input_data[201]
  PIN input_data[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 665.250 796.000 665.530 800.000 ;
    END
  END input_data[202]
  PIN input_data[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 668.470 796.000 668.750 800.000 ;
    END
  END input_data[203]
  PIN input_data[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 671.690 796.000 671.970 800.000 ;
    END
  END input_data[204]
  PIN input_data[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 674.910 796.000 675.190 800.000 ;
    END
  END input_data[205]
  PIN input_data[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 678.130 796.000 678.410 800.000 ;
    END
  END input_data[206]
  PIN input_data[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 681.350 796.000 681.630 800.000 ;
    END
  END input_data[207]
  PIN input_data[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 684.570 796.000 684.850 800.000 ;
    END
  END input_data[208]
  PIN input_data[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 687.790 796.000 688.070 800.000 ;
    END
  END input_data[209]
  PIN input_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 79.210 796.000 79.490 800.000 ;
    END
  END input_data[20]
  PIN input_data[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 691.010 796.000 691.290 800.000 ;
    END
  END input_data[210]
  PIN input_data[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 694.230 796.000 694.510 800.000 ;
    END
  END input_data[211]
  PIN input_data[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 697.450 796.000 697.730 800.000 ;
    END
  END input_data[212]
  PIN input_data[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 700.670 796.000 700.950 800.000 ;
    END
  END input_data[213]
  PIN input_data[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 703.890 796.000 704.170 800.000 ;
    END
  END input_data[214]
  PIN input_data[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 707.110 796.000 707.390 800.000 ;
    END
  END input_data[215]
  PIN input_data[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 710.330 796.000 710.610 800.000 ;
    END
  END input_data[216]
  PIN input_data[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 713.550 796.000 713.830 800.000 ;
    END
  END input_data[217]
  PIN input_data[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 716.770 796.000 717.050 800.000 ;
    END
  END input_data[218]
  PIN input_data[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 719.990 796.000 720.270 800.000 ;
    END
  END input_data[219]
  PIN input_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.430 796.000 82.710 800.000 ;
    END
  END input_data[21]
  PIN input_data[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 723.210 796.000 723.490 800.000 ;
    END
  END input_data[220]
  PIN input_data[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 726.430 796.000 726.710 800.000 ;
    END
  END input_data[221]
  PIN input_data[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 729.650 796.000 729.930 800.000 ;
    END
  END input_data[222]
  PIN input_data[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 796.000 733.150 800.000 ;
    END
  END input_data[223]
  PIN input_data[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 736.090 796.000 736.370 800.000 ;
    END
  END input_data[224]
  PIN input_data[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 739.310 796.000 739.590 800.000 ;
    END
  END input_data[225]
  PIN input_data[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 742.530 796.000 742.810 800.000 ;
    END
  END input_data[226]
  PIN input_data[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 745.750 796.000 746.030 800.000 ;
    END
  END input_data[227]
  PIN input_data[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 748.970 796.000 749.250 800.000 ;
    END
  END input_data[228]
  PIN input_data[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 752.190 796.000 752.470 800.000 ;
    END
  END input_data[229]
  PIN input_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.650 796.000 85.930 800.000 ;
    END
  END input_data[22]
  PIN input_data[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 755.410 796.000 755.690 800.000 ;
    END
  END input_data[230]
  PIN input_data[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 758.630 796.000 758.910 800.000 ;
    END
  END input_data[231]
  PIN input_data[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 761.850 796.000 762.130 800.000 ;
    END
  END input_data[232]
  PIN input_data[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 765.070 796.000 765.350 800.000 ;
    END
  END input_data[233]
  PIN input_data[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 768.290 796.000 768.570 800.000 ;
    END
  END input_data[234]
  PIN input_data[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 771.510 796.000 771.790 800.000 ;
    END
  END input_data[235]
  PIN input_data[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 774.730 796.000 775.010 800.000 ;
    END
  END input_data[236]
  PIN input_data[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 777.950 796.000 778.230 800.000 ;
    END
  END input_data[237]
  PIN input_data[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 796.000 781.450 800.000 ;
    END
  END input_data[238]
  PIN input_data[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 796.000 784.670 800.000 ;
    END
  END input_data[239]
  PIN input_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.870 796.000 89.150 800.000 ;
    END
  END input_data[23]
  PIN input_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 92.090 796.000 92.370 800.000 ;
    END
  END input_data[24]
  PIN input_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 95.310 796.000 95.590 800.000 ;
    END
  END input_data[25]
  PIN input_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 98.530 796.000 98.810 800.000 ;
    END
  END input_data[26]
  PIN input_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 101.750 796.000 102.030 800.000 ;
    END
  END input_data[27]
  PIN input_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 104.970 796.000 105.250 800.000 ;
    END
  END input_data[28]
  PIN input_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 108.190 796.000 108.470 800.000 ;
    END
  END input_data[29]
  PIN input_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 21.250 796.000 21.530 800.000 ;
    END
  END input_data[2]
  PIN input_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 111.410 796.000 111.690 800.000 ;
    END
  END input_data[30]
  PIN input_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 114.630 796.000 114.910 800.000 ;
    END
  END input_data[31]
  PIN input_data[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 117.850 796.000 118.130 800.000 ;
    END
  END input_data[32]
  PIN input_data[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 121.070 796.000 121.350 800.000 ;
    END
  END input_data[33]
  PIN input_data[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.290 796.000 124.570 800.000 ;
    END
  END input_data[34]
  PIN input_data[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 127.510 796.000 127.790 800.000 ;
    END
  END input_data[35]
  PIN input_data[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 130.730 796.000 131.010 800.000 ;
    END
  END input_data[36]
  PIN input_data[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 133.950 796.000 134.230 800.000 ;
    END
  END input_data[37]
  PIN input_data[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 137.170 796.000 137.450 800.000 ;
    END
  END input_data[38]
  PIN input_data[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.390 796.000 140.670 800.000 ;
    END
  END input_data[39]
  PIN input_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 24.470 796.000 24.750 800.000 ;
    END
  END input_data[3]
  PIN input_data[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 143.610 796.000 143.890 800.000 ;
    END
  END input_data[40]
  PIN input_data[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 146.830 796.000 147.110 800.000 ;
    END
  END input_data[41]
  PIN input_data[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 150.050 796.000 150.330 800.000 ;
    END
  END input_data[42]
  PIN input_data[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 153.270 796.000 153.550 800.000 ;
    END
  END input_data[43]
  PIN input_data[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 156.490 796.000 156.770 800.000 ;
    END
  END input_data[44]
  PIN input_data[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 159.710 796.000 159.990 800.000 ;
    END
  END input_data[45]
  PIN input_data[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.930 796.000 163.210 800.000 ;
    END
  END input_data[46]
  PIN input_data[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 166.150 796.000 166.430 800.000 ;
    END
  END input_data[47]
  PIN input_data[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.370 796.000 169.650 800.000 ;
    END
  END input_data[48]
  PIN input_data[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 172.590 796.000 172.870 800.000 ;
    END
  END input_data[49]
  PIN input_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 27.690 796.000 27.970 800.000 ;
    END
  END input_data[4]
  PIN input_data[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.810 796.000 176.090 800.000 ;
    END
  END input_data[50]
  PIN input_data[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 179.030 796.000 179.310 800.000 ;
    END
  END input_data[51]
  PIN input_data[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 182.250 796.000 182.530 800.000 ;
    END
  END input_data[52]
  PIN input_data[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 185.470 796.000 185.750 800.000 ;
    END
  END input_data[53]
  PIN input_data[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 188.690 796.000 188.970 800.000 ;
    END
  END input_data[54]
  PIN input_data[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.910 796.000 192.190 800.000 ;
    END
  END input_data[55]
  PIN input_data[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.130 796.000 195.410 800.000 ;
    END
  END input_data[56]
  PIN input_data[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 198.350 796.000 198.630 800.000 ;
    END
  END input_data[57]
  PIN input_data[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 201.570 796.000 201.850 800.000 ;
    END
  END input_data[58]
  PIN input_data[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 204.790 796.000 205.070 800.000 ;
    END
  END input_data[59]
  PIN input_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 30.910 796.000 31.190 800.000 ;
    END
  END input_data[5]
  PIN input_data[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 208.010 796.000 208.290 800.000 ;
    END
  END input_data[60]
  PIN input_data[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 211.230 796.000 211.510 800.000 ;
    END
  END input_data[61]
  PIN input_data[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 214.450 796.000 214.730 800.000 ;
    END
  END input_data[62]
  PIN input_data[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.670 796.000 217.950 800.000 ;
    END
  END input_data[63]
  PIN input_data[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 220.890 796.000 221.170 800.000 ;
    END
  END input_data[64]
  PIN input_data[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 224.110 796.000 224.390 800.000 ;
    END
  END input_data[65]
  PIN input_data[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 227.330 796.000 227.610 800.000 ;
    END
  END input_data[66]
  PIN input_data[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 230.550 796.000 230.830 800.000 ;
    END
  END input_data[67]
  PIN input_data[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 233.770 796.000 234.050 800.000 ;
    END
  END input_data[68]
  PIN input_data[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 236.990 796.000 237.270 800.000 ;
    END
  END input_data[69]
  PIN input_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 34.130 796.000 34.410 800.000 ;
    END
  END input_data[6]
  PIN input_data[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 240.210 796.000 240.490 800.000 ;
    END
  END input_data[70]
  PIN input_data[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 243.430 796.000 243.710 800.000 ;
    END
  END input_data[71]
  PIN input_data[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 246.650 796.000 246.930 800.000 ;
    END
  END input_data[72]
  PIN input_data[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 249.870 796.000 250.150 800.000 ;
    END
  END input_data[73]
  PIN input_data[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 253.090 796.000 253.370 800.000 ;
    END
  END input_data[74]
  PIN input_data[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 256.310 796.000 256.590 800.000 ;
    END
  END input_data[75]
  PIN input_data[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 259.530 796.000 259.810 800.000 ;
    END
  END input_data[76]
  PIN input_data[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 262.750 796.000 263.030 800.000 ;
    END
  END input_data[77]
  PIN input_data[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 265.970 796.000 266.250 800.000 ;
    END
  END input_data[78]
  PIN input_data[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 269.190 796.000 269.470 800.000 ;
    END
  END input_data[79]
  PIN input_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 37.350 796.000 37.630 800.000 ;
    END
  END input_data[7]
  PIN input_data[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 272.410 796.000 272.690 800.000 ;
    END
  END input_data[80]
  PIN input_data[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 275.630 796.000 275.910 800.000 ;
    END
  END input_data[81]
  PIN input_data[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 278.850 796.000 279.130 800.000 ;
    END
  END input_data[82]
  PIN input_data[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 282.070 796.000 282.350 800.000 ;
    END
  END input_data[83]
  PIN input_data[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 285.290 796.000 285.570 800.000 ;
    END
  END input_data[84]
  PIN input_data[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 288.510 796.000 288.790 800.000 ;
    END
  END input_data[85]
  PIN input_data[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 291.730 796.000 292.010 800.000 ;
    END
  END input_data[86]
  PIN input_data[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 294.950 796.000 295.230 800.000 ;
    END
  END input_data[87]
  PIN input_data[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 298.170 796.000 298.450 800.000 ;
    END
  END input_data[88]
  PIN input_data[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 301.390 796.000 301.670 800.000 ;
    END
  END input_data[89]
  PIN input_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 40.570 796.000 40.850 800.000 ;
    END
  END input_data[8]
  PIN input_data[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 304.610 796.000 304.890 800.000 ;
    END
  END input_data[90]
  PIN input_data[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 307.830 796.000 308.110 800.000 ;
    END
  END input_data[91]
  PIN input_data[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 311.050 796.000 311.330 800.000 ;
    END
  END input_data[92]
  PIN input_data[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 314.270 796.000 314.550 800.000 ;
    END
  END input_data[93]
  PIN input_data[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 317.490 796.000 317.770 800.000 ;
    END
  END input_data[94]
  PIN input_data[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 320.710 796.000 320.990 800.000 ;
    END
  END input_data[95]
  PIN input_data[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 323.930 796.000 324.210 800.000 ;
    END
  END input_data[96]
  PIN input_data[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 327.150 796.000 327.430 800.000 ;
    END
  END input_data[97]
  PIN input_data[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 330.370 796.000 330.650 800.000 ;
    END
  END input_data[98]
  PIN input_data[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 333.590 796.000 333.870 800.000 ;
    END
  END input_data[99]
  PIN input_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 43.790 796.000 44.070 800.000 ;
    END
  END input_data[9]
  PIN output_low[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END output_low[0]
  PIN output_low[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END output_low[10]
  PIN output_low[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END output_low[11]
  PIN output_low[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END output_low[12]
  PIN output_low[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END output_low[13]
  PIN output_low[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END output_low[14]
  PIN output_low[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END output_low[15]
  PIN output_low[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END output_low[1]
  PIN output_low[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END output_low[2]
  PIN output_low[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END output_low[3]
  PIN output_low[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END output_low[4]
  PIN output_low[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END output_low[5]
  PIN output_low[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END output_low[6]
  PIN output_low[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END output_low[7]
  PIN output_low[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.000 4.000 423.600 ;
    END
  END output_low[8]
  PIN output_low[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.960 4.000 472.560 ;
    END
  END output_low[9]
  PIN tap[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END tap[0]
  PIN tap[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END tap[1]
  PIN tap[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END tap[2]
  PIN tap[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END tap[3]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 788.885 ;
      LAYER met1 ;
        RECT 3.750 10.640 794.720 790.460 ;
      LAYER met2 ;
        RECT 3.770 795.720 14.530 796.690 ;
        RECT 15.370 795.720 17.750 796.690 ;
        RECT 18.590 795.720 20.970 796.690 ;
        RECT 21.810 795.720 24.190 796.690 ;
        RECT 25.030 795.720 27.410 796.690 ;
        RECT 28.250 795.720 30.630 796.690 ;
        RECT 31.470 795.720 33.850 796.690 ;
        RECT 34.690 795.720 37.070 796.690 ;
        RECT 37.910 795.720 40.290 796.690 ;
        RECT 41.130 795.720 43.510 796.690 ;
        RECT 44.350 795.720 46.730 796.690 ;
        RECT 47.570 795.720 49.950 796.690 ;
        RECT 50.790 795.720 53.170 796.690 ;
        RECT 54.010 795.720 56.390 796.690 ;
        RECT 57.230 795.720 59.610 796.690 ;
        RECT 60.450 795.720 62.830 796.690 ;
        RECT 63.670 795.720 66.050 796.690 ;
        RECT 66.890 795.720 69.270 796.690 ;
        RECT 70.110 795.720 72.490 796.690 ;
        RECT 73.330 795.720 75.710 796.690 ;
        RECT 76.550 795.720 78.930 796.690 ;
        RECT 79.770 795.720 82.150 796.690 ;
        RECT 82.990 795.720 85.370 796.690 ;
        RECT 86.210 795.720 88.590 796.690 ;
        RECT 89.430 795.720 91.810 796.690 ;
        RECT 92.650 795.720 95.030 796.690 ;
        RECT 95.870 795.720 98.250 796.690 ;
        RECT 99.090 795.720 101.470 796.690 ;
        RECT 102.310 795.720 104.690 796.690 ;
        RECT 105.530 795.720 107.910 796.690 ;
        RECT 108.750 795.720 111.130 796.690 ;
        RECT 111.970 795.720 114.350 796.690 ;
        RECT 115.190 795.720 117.570 796.690 ;
        RECT 118.410 795.720 120.790 796.690 ;
        RECT 121.630 795.720 124.010 796.690 ;
        RECT 124.850 795.720 127.230 796.690 ;
        RECT 128.070 795.720 130.450 796.690 ;
        RECT 131.290 795.720 133.670 796.690 ;
        RECT 134.510 795.720 136.890 796.690 ;
        RECT 137.730 795.720 140.110 796.690 ;
        RECT 140.950 795.720 143.330 796.690 ;
        RECT 144.170 795.720 146.550 796.690 ;
        RECT 147.390 795.720 149.770 796.690 ;
        RECT 150.610 795.720 152.990 796.690 ;
        RECT 153.830 795.720 156.210 796.690 ;
        RECT 157.050 795.720 159.430 796.690 ;
        RECT 160.270 795.720 162.650 796.690 ;
        RECT 163.490 795.720 165.870 796.690 ;
        RECT 166.710 795.720 169.090 796.690 ;
        RECT 169.930 795.720 172.310 796.690 ;
        RECT 173.150 795.720 175.530 796.690 ;
        RECT 176.370 795.720 178.750 796.690 ;
        RECT 179.590 795.720 181.970 796.690 ;
        RECT 182.810 795.720 185.190 796.690 ;
        RECT 186.030 795.720 188.410 796.690 ;
        RECT 189.250 795.720 191.630 796.690 ;
        RECT 192.470 795.720 194.850 796.690 ;
        RECT 195.690 795.720 198.070 796.690 ;
        RECT 198.910 795.720 201.290 796.690 ;
        RECT 202.130 795.720 204.510 796.690 ;
        RECT 205.350 795.720 207.730 796.690 ;
        RECT 208.570 795.720 210.950 796.690 ;
        RECT 211.790 795.720 214.170 796.690 ;
        RECT 215.010 795.720 217.390 796.690 ;
        RECT 218.230 795.720 220.610 796.690 ;
        RECT 221.450 795.720 223.830 796.690 ;
        RECT 224.670 795.720 227.050 796.690 ;
        RECT 227.890 795.720 230.270 796.690 ;
        RECT 231.110 795.720 233.490 796.690 ;
        RECT 234.330 795.720 236.710 796.690 ;
        RECT 237.550 795.720 239.930 796.690 ;
        RECT 240.770 795.720 243.150 796.690 ;
        RECT 243.990 795.720 246.370 796.690 ;
        RECT 247.210 795.720 249.590 796.690 ;
        RECT 250.430 795.720 252.810 796.690 ;
        RECT 253.650 795.720 256.030 796.690 ;
        RECT 256.870 795.720 259.250 796.690 ;
        RECT 260.090 795.720 262.470 796.690 ;
        RECT 263.310 795.720 265.690 796.690 ;
        RECT 266.530 795.720 268.910 796.690 ;
        RECT 269.750 795.720 272.130 796.690 ;
        RECT 272.970 795.720 275.350 796.690 ;
        RECT 276.190 795.720 278.570 796.690 ;
        RECT 279.410 795.720 281.790 796.690 ;
        RECT 282.630 795.720 285.010 796.690 ;
        RECT 285.850 795.720 288.230 796.690 ;
        RECT 289.070 795.720 291.450 796.690 ;
        RECT 292.290 795.720 294.670 796.690 ;
        RECT 295.510 795.720 297.890 796.690 ;
        RECT 298.730 795.720 301.110 796.690 ;
        RECT 301.950 795.720 304.330 796.690 ;
        RECT 305.170 795.720 307.550 796.690 ;
        RECT 308.390 795.720 310.770 796.690 ;
        RECT 311.610 795.720 313.990 796.690 ;
        RECT 314.830 795.720 317.210 796.690 ;
        RECT 318.050 795.720 320.430 796.690 ;
        RECT 321.270 795.720 323.650 796.690 ;
        RECT 324.490 795.720 326.870 796.690 ;
        RECT 327.710 795.720 330.090 796.690 ;
        RECT 330.930 795.720 333.310 796.690 ;
        RECT 334.150 795.720 336.530 796.690 ;
        RECT 337.370 795.720 339.750 796.690 ;
        RECT 340.590 795.720 342.970 796.690 ;
        RECT 343.810 795.720 346.190 796.690 ;
        RECT 347.030 795.720 349.410 796.690 ;
        RECT 350.250 795.720 352.630 796.690 ;
        RECT 353.470 795.720 355.850 796.690 ;
        RECT 356.690 795.720 359.070 796.690 ;
        RECT 359.910 795.720 362.290 796.690 ;
        RECT 363.130 795.720 365.510 796.690 ;
        RECT 366.350 795.720 368.730 796.690 ;
        RECT 369.570 795.720 371.950 796.690 ;
        RECT 372.790 795.720 375.170 796.690 ;
        RECT 376.010 795.720 378.390 796.690 ;
        RECT 379.230 795.720 381.610 796.690 ;
        RECT 382.450 795.720 384.830 796.690 ;
        RECT 385.670 795.720 388.050 796.690 ;
        RECT 388.890 795.720 391.270 796.690 ;
        RECT 392.110 795.720 394.490 796.690 ;
        RECT 395.330 795.720 397.710 796.690 ;
        RECT 398.550 795.720 400.930 796.690 ;
        RECT 401.770 795.720 404.150 796.690 ;
        RECT 404.990 795.720 407.370 796.690 ;
        RECT 408.210 795.720 410.590 796.690 ;
        RECT 411.430 795.720 413.810 796.690 ;
        RECT 414.650 795.720 417.030 796.690 ;
        RECT 417.870 795.720 420.250 796.690 ;
        RECT 421.090 795.720 423.470 796.690 ;
        RECT 424.310 795.720 426.690 796.690 ;
        RECT 427.530 795.720 429.910 796.690 ;
        RECT 430.750 795.720 433.130 796.690 ;
        RECT 433.970 795.720 436.350 796.690 ;
        RECT 437.190 795.720 439.570 796.690 ;
        RECT 440.410 795.720 442.790 796.690 ;
        RECT 443.630 795.720 446.010 796.690 ;
        RECT 446.850 795.720 449.230 796.690 ;
        RECT 450.070 795.720 452.450 796.690 ;
        RECT 453.290 795.720 455.670 796.690 ;
        RECT 456.510 795.720 458.890 796.690 ;
        RECT 459.730 795.720 462.110 796.690 ;
        RECT 462.950 795.720 465.330 796.690 ;
        RECT 466.170 795.720 468.550 796.690 ;
        RECT 469.390 795.720 471.770 796.690 ;
        RECT 472.610 795.720 474.990 796.690 ;
        RECT 475.830 795.720 478.210 796.690 ;
        RECT 479.050 795.720 481.430 796.690 ;
        RECT 482.270 795.720 484.650 796.690 ;
        RECT 485.490 795.720 487.870 796.690 ;
        RECT 488.710 795.720 491.090 796.690 ;
        RECT 491.930 795.720 494.310 796.690 ;
        RECT 495.150 795.720 497.530 796.690 ;
        RECT 498.370 795.720 500.750 796.690 ;
        RECT 501.590 795.720 503.970 796.690 ;
        RECT 504.810 795.720 507.190 796.690 ;
        RECT 508.030 795.720 510.410 796.690 ;
        RECT 511.250 795.720 513.630 796.690 ;
        RECT 514.470 795.720 516.850 796.690 ;
        RECT 517.690 795.720 520.070 796.690 ;
        RECT 520.910 795.720 523.290 796.690 ;
        RECT 524.130 795.720 526.510 796.690 ;
        RECT 527.350 795.720 529.730 796.690 ;
        RECT 530.570 795.720 532.950 796.690 ;
        RECT 533.790 795.720 536.170 796.690 ;
        RECT 537.010 795.720 539.390 796.690 ;
        RECT 540.230 795.720 542.610 796.690 ;
        RECT 543.450 795.720 545.830 796.690 ;
        RECT 546.670 795.720 549.050 796.690 ;
        RECT 549.890 795.720 552.270 796.690 ;
        RECT 553.110 795.720 555.490 796.690 ;
        RECT 556.330 795.720 558.710 796.690 ;
        RECT 559.550 795.720 561.930 796.690 ;
        RECT 562.770 795.720 565.150 796.690 ;
        RECT 565.990 795.720 568.370 796.690 ;
        RECT 569.210 795.720 571.590 796.690 ;
        RECT 572.430 795.720 574.810 796.690 ;
        RECT 575.650 795.720 578.030 796.690 ;
        RECT 578.870 795.720 581.250 796.690 ;
        RECT 582.090 795.720 584.470 796.690 ;
        RECT 585.310 795.720 587.690 796.690 ;
        RECT 588.530 795.720 590.910 796.690 ;
        RECT 591.750 795.720 594.130 796.690 ;
        RECT 594.970 795.720 597.350 796.690 ;
        RECT 598.190 795.720 600.570 796.690 ;
        RECT 601.410 795.720 603.790 796.690 ;
        RECT 604.630 795.720 607.010 796.690 ;
        RECT 607.850 795.720 610.230 796.690 ;
        RECT 611.070 795.720 613.450 796.690 ;
        RECT 614.290 795.720 616.670 796.690 ;
        RECT 617.510 795.720 619.890 796.690 ;
        RECT 620.730 795.720 623.110 796.690 ;
        RECT 623.950 795.720 626.330 796.690 ;
        RECT 627.170 795.720 629.550 796.690 ;
        RECT 630.390 795.720 632.770 796.690 ;
        RECT 633.610 795.720 635.990 796.690 ;
        RECT 636.830 795.720 639.210 796.690 ;
        RECT 640.050 795.720 642.430 796.690 ;
        RECT 643.270 795.720 645.650 796.690 ;
        RECT 646.490 795.720 648.870 796.690 ;
        RECT 649.710 795.720 652.090 796.690 ;
        RECT 652.930 795.720 655.310 796.690 ;
        RECT 656.150 795.720 658.530 796.690 ;
        RECT 659.370 795.720 661.750 796.690 ;
        RECT 662.590 795.720 664.970 796.690 ;
        RECT 665.810 795.720 668.190 796.690 ;
        RECT 669.030 795.720 671.410 796.690 ;
        RECT 672.250 795.720 674.630 796.690 ;
        RECT 675.470 795.720 677.850 796.690 ;
        RECT 678.690 795.720 681.070 796.690 ;
        RECT 681.910 795.720 684.290 796.690 ;
        RECT 685.130 795.720 687.510 796.690 ;
        RECT 688.350 795.720 690.730 796.690 ;
        RECT 691.570 795.720 693.950 796.690 ;
        RECT 694.790 795.720 697.170 796.690 ;
        RECT 698.010 795.720 700.390 796.690 ;
        RECT 701.230 795.720 703.610 796.690 ;
        RECT 704.450 795.720 706.830 796.690 ;
        RECT 707.670 795.720 710.050 796.690 ;
        RECT 710.890 795.720 713.270 796.690 ;
        RECT 714.110 795.720 716.490 796.690 ;
        RECT 717.330 795.720 719.710 796.690 ;
        RECT 720.550 795.720 722.930 796.690 ;
        RECT 723.770 795.720 726.150 796.690 ;
        RECT 726.990 795.720 729.370 796.690 ;
        RECT 730.210 795.720 732.590 796.690 ;
        RECT 733.430 795.720 735.810 796.690 ;
        RECT 736.650 795.720 739.030 796.690 ;
        RECT 739.870 795.720 742.250 796.690 ;
        RECT 743.090 795.720 745.470 796.690 ;
        RECT 746.310 795.720 748.690 796.690 ;
        RECT 749.530 795.720 751.910 796.690 ;
        RECT 752.750 795.720 755.130 796.690 ;
        RECT 755.970 795.720 758.350 796.690 ;
        RECT 759.190 795.720 761.570 796.690 ;
        RECT 762.410 795.720 764.790 796.690 ;
        RECT 765.630 795.720 768.010 796.690 ;
        RECT 768.850 795.720 771.230 796.690 ;
        RECT 772.070 795.720 774.450 796.690 ;
        RECT 775.290 795.720 777.670 796.690 ;
        RECT 778.510 795.720 780.890 796.690 ;
        RECT 781.730 795.720 784.110 796.690 ;
        RECT 784.950 795.720 793.910 796.690 ;
        RECT 3.770 4.280 793.910 795.720 ;
        RECT 3.770 4.000 100.090 4.280 ;
        RECT 100.930 4.000 299.730 4.280 ;
        RECT 300.570 4.000 499.370 4.280 ;
        RECT 500.210 4.000 699.010 4.280 ;
        RECT 699.850 4.000 793.910 4.280 ;
      LAYER met3 ;
        RECT 3.745 766.720 796.000 788.965 ;
        RECT 4.400 765.320 796.000 766.720 ;
        RECT 3.745 717.760 796.000 765.320 ;
        RECT 4.400 716.360 796.000 717.760 ;
        RECT 3.745 668.800 796.000 716.360 ;
        RECT 4.400 667.400 796.000 668.800 ;
        RECT 3.745 619.840 796.000 667.400 ;
        RECT 4.400 618.440 796.000 619.840 ;
        RECT 3.745 570.880 796.000 618.440 ;
        RECT 4.400 569.480 796.000 570.880 ;
        RECT 3.745 521.920 796.000 569.480 ;
        RECT 4.400 520.520 796.000 521.920 ;
        RECT 3.745 472.960 796.000 520.520 ;
        RECT 4.400 471.560 796.000 472.960 ;
        RECT 3.745 424.000 796.000 471.560 ;
        RECT 4.400 422.600 796.000 424.000 ;
        RECT 3.745 399.520 796.000 422.600 ;
        RECT 3.745 398.120 795.600 399.520 ;
        RECT 3.745 375.040 796.000 398.120 ;
        RECT 4.400 373.640 796.000 375.040 ;
        RECT 3.745 326.080 796.000 373.640 ;
        RECT 4.400 324.680 796.000 326.080 ;
        RECT 3.745 277.120 796.000 324.680 ;
        RECT 4.400 275.720 796.000 277.120 ;
        RECT 3.745 228.160 796.000 275.720 ;
        RECT 4.400 226.760 796.000 228.160 ;
        RECT 3.745 179.200 796.000 226.760 ;
        RECT 4.400 177.800 796.000 179.200 ;
        RECT 3.745 130.240 796.000 177.800 ;
        RECT 4.400 128.840 796.000 130.240 ;
        RECT 3.745 81.280 796.000 128.840 ;
        RECT 4.400 79.880 796.000 81.280 ;
        RECT 3.745 32.320 796.000 79.880 ;
        RECT 4.400 30.920 796.000 32.320 ;
        RECT 3.745 10.715 796.000 30.920 ;
      LAYER met4 ;
        RECT 3.975 136.855 20.640 787.945 ;
        RECT 23.040 136.855 23.940 787.945 ;
        RECT 26.340 136.855 174.240 787.945 ;
        RECT 176.640 136.855 177.540 787.945 ;
        RECT 179.940 136.855 327.840 787.945 ;
        RECT 330.240 136.855 331.140 787.945 ;
        RECT 333.540 136.855 481.440 787.945 ;
        RECT 483.840 136.855 484.740 787.945 ;
        RECT 487.140 136.855 635.040 787.945 ;
        RECT 637.440 136.855 638.340 787.945 ;
        RECT 640.740 136.855 743.065 787.945 ;
  END
END lowpass
END LIBRARY

